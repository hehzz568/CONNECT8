// vga_controller.v — 8x8 to 640x480
module vga_controller(
    input  wire        clk, reset,
    input  wire [63:0] game_grid,
    input  wire [63:0] block1, block2, block3,
    input  wire [2:0]  block1_x, block1_y,
    input  wire [2:0]  block2_x, block2_y,
    input  wire [2:0]  block3_x, block3_y,
    input  wire [7:0]  score,
    input  wire        game_over,
    input  wire        show_title,         
    output reg  [7:0]  vga_r, vga_g, vga_b,
    output wire        vga_hs, vga_vs, vga_blank_n
);
    wire [9:0] x, y;
    vga_timing_640x480 T(
        .clk(clk), .reset(reset),
        .x(x), .y(y),
        .hs(vga_hs), .vs(vga_vs), .blank_n(vga_blank_n)
    );

    // title ROM (splash image) 
    wire [18:0] title_addr = y * 10'd640 + x;
    wire [7:0]  title_idx;

    // IP generated by MegaWizard: title_rom
    title_rom U_TITLE (
        .address(title_addr),
        .clock  (clk),
        .q      (title_idx)
    );

    // simple palette: index -> RGB
    reg [7:0] title_r, title_g, title_b;
    always @* begin
        case (title_idx)
            8'd0: begin            // dark blue background
                title_r = 8'd15;
                title_g = 8'd45;
                title_b = 8'd82;
            end
            8'd1: begin            // light yellow panel
                title_r = 8'd217;
                title_g = 8'd201;
                title_b = 8'd143;
            end
            8'd2: begin            // blue text
                title_r = 8'd27;
                title_g = 8'd78;
                title_b = 8'd142;
            end
            default: begin
                title_r = 8'd0;
                title_g = 8'd0;
                title_b = 8'd0;
            end
        endcase
    end

    // 8x8, each 80x60
    wire [2:0] cell_x = x/80;
    wire [2:0] cell_y = y/60;
    wire [6:0] idx    = cell_y*8 + cell_x;

    // block on line
    wire on_vline = (x%80==0);
    wire on_hline = (y%60==0);
    wire on_grid  = on_vline || on_hline;

    // shadow for these 3
    function inside_block;
        input [63:0] blk; input [2:0] bx, by; input [2:0] cx, cy;
        integer i,j;
        reg hit;
        begin
            hit = 0;
            for (i=0;i<8;i=i+1) begin
                for (j=0;j<8;j=j+1) begin
                    if (blk[i*8+j]) begin
                        if ((bx+j)==cx && (by+i)==cy) hit=1;
                    end
                end
            end
            inside_block = hit;
        end
    endfunction

    wire grid_on = game_grid[idx];
    wire blk1_on = inside_block(block1,block1_x,block1_y,cell_x,cell_y);
    wire blk2_on = inside_block(block2,block2_x,block2_y,cell_x,cell_y);
    wire blk3_on = inside_block(block3,block3_x,block3_y,cell_x,cell_y);

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            vga_r <= 0; vga_g <= 0; vga_b <= 0;
        end
        else if (!vga_blank_n) begin
            vga_r <= 0; vga_g <= 0; vga_b <= 0;
        end
        else begin
            if (show_title) begin
                // show splash image
                vga_r <= title_r;
                vga_g <= title_g;
                vga_b <= title_b;
            end
            else if (grid_on) begin
                {vga_r,vga_g,vga_b} <= {8'hE0,8'h60,8'h20}; // placed: orange
            end
            else if (blk1_on|blk2_on|blk3_on) begin
                {vga_r,vga_g,vga_b} <= {8'h80,8'hC0,8'hFF}; // pending: blue
            end
            else if (on_grid) begin
                {vga_r,vga_g,vga_b} <= {8'h40,8'h40,8'h40}; // line: grey
            end
            else begin
                {vga_r,vga_g,vga_b} <= 24'h000000;          // background: black
            end
        end
    end
endmodule

